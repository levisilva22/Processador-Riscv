//COMPILE: iverilog.exe -g2012 -o riscvsingle_p1.vcd -tvvp .\riscvsingle_p1.sv
//SIMULATE: vvp riscvsingle_p1

// Implementa toda a arquitetura do riscv
module top(input  logic        clk, reset, 
           output logic [31:0] WriteData, DataAdr, 
           output logic        MemWrite);

  logic [31:0] PC, Instr, ReadData;
  
  // instantiate processor and memories
  riscvsingle rvsingle(clk, reset, PC, Instr, MemWrite, DataAdr, 
                       WriteData, ReadData);
  imem imem(PC, Instr); // instancia a memória de instrução
  dmem dmem(clk, MemWrite, DataAdr, WriteData, ReadData); // instancia a memória de dados
endmodule

module riscvsingle(input  logic        clk, reset,
                   output logic [31:0] PC,
                   input  logic [31:0] Instr,
                   output logic        MemWrite,
                   output logic [31:0] ALUResult, WriteData,
                   input  logic [31:0] ReadData);
  // sinal do bloco de controle
  logic       ALUSrc, RegWrite, Jump, Zero;
  logic [1:0] ResultSrc, ImmSrc;
  logic [2:0] ALUControl;

  controller c(Instr[6:0], Instr[14:12], Instr[30], Zero,
               ResultSrc, MemWrite, PCSrc,
               ALUSrc, RegWrite, Jump,
               ImmSrc, ALUControl); // Gera os sinal de controle 
  datapath dp(clk, reset, ResultSrc, PCSrc,
              ALUSrc, RegWrite,
              ImmSrc, ALUControl,
              Zero, PC, Instr,
              ALUResult, WriteData, ReadData);
endmodule

// Modulo para gerar os sinal de controle
module controller(input  logic [6:0] op,
                  input  logic [2:0] funct3,
                  input  logic       funct7b5,
                  input  logic       Zero,
                  output logic [1:0] ResultSrc,
                  output logic       MemWrite,
                  output logic       PCSrc, ALUSrc,
                  output logic       RegWrite, Jump,
                  output logic [1:0] ImmSrc,
                  output logic [2:0] ALUControl);

  logic [1:0] ALUOp;
  logic       Branch;
  
  /* 
    A função do bloco de controle é decodificar os bits da instrução
    com isso maindec e aludec decoficam qual será a instrução e qual operação será feita 
    na ALU, respectivamente
  */
  maindec md(op, ResultSrc, MemWrite, Branch,
             ALUSrc, RegWrite, Jump, ImmSrc, ALUOp); //decodifica a operação a ser realizada
  aludec  ad(op[5], funct3, funct7b5, ALUOp, ALUControl);

  assign PCSrc = Branch & Zero; // PCsrc só ocorre se branch e a operação de subtração na ALU for zero
endmodule

// Modulo para decodificar a instrução
module maindec(input  logic [6:0] op,
               output logic [1:0] ResultSrc,
               output logic       MemWrite,
               output logic       Branch, ALUSrc,
               output logic       RegWrite, Jump,
               output logic [1:0] ImmSrc,
               output logic [1:0] ALUOp);

  logic [11:0] controls; // instancia um array de 11 bits 

  assign {RegWrite, ImmSrc, ALUSrc, MemWrite,
          ResultSrc, Branch, ALUOp, Jump} = controls; //atribui os bits recebido ao controle 

  always_comb 
    case(op)
    // RegWrite_ImmSrc_ALUSrc_MemWrite_ResultSrc_Branch_ALUOp_Jump
      7'b0000011: controls = 12'b1_00_1_0_01_0_00_0; // lw
      7'b0100011: controls = 12'b0_01_1_1_00_0_00_0; // sw
      7'b0110011: controls = 12'b1_xx_0_0_00_0_10_0; // R-type
      7'b1100011: controls = 12'b0_10_0_0_00_1_01_0; // beq
      7'b0010011: controls = 12'b1_00_1_0_00_0_10_0; // I-type ALU (addi, etc.)
      7'b1101111: controls = 12'b1_11_0_0_10_0_00_1; // jal
      default:    controls = 12'bx_xx_x_x_xx_x_xx_x; // non-implemented instruction
    endcase
endmodule

// modulo de decodifica a operação feita na alu
module aludec(input  logic       opb5,
              input  logic [2:0] funct3,
              input  logic       funct7b5, 
              input  logic [1:0] ALUOp,
              output logic [2:0] ALUControl);

  logic  RtypeSub;
  // se o 5 bit dos 7 bits de funct7 for 1 e se o bit 5 de opcode for 1
  assign RtypeSub = funct7b5 & opb5;  // TRUE for R-type subtract instruction

  always_comb
    case(ALUOp)
      2'b00:                ALUControl = 3'b000; // addition, lw, sw
      2'b01:                ALUControl = 3'b001; // subtraction, branch
      default: case(funct3) // R-type or I-type ALU
                 3'b000:  if (RtypeSub) 
                            ALUControl = 3'b001; // sub
                          else          
                            ALUControl = 3'b000; // add, addi
                 3'b010:    ALUControl = 3'b101; // slt, slti
                 3'b110:    ALUControl = 3'b011; // or, ori
                 3'b111:    ALUControl = 3'b010; // and, andi
                 default:   ALUControl = 3'bxxx; // ???
               endcase
    endcase
endmodule

module datapath(input  logic        clk, reset,
                input  logic [1:0]  ResultSrc, 
                input  logic        PCSrc, ALUSrc,
                input  logic        RegWrite,
                input  logic [1:0]  ImmSrc,
                input  logic [2:0]  ALUControl,
                output logic        Zero,
                output logic [31:0] PC,
                input  logic [31:0] Instr,
                output logic [31:0] ALUResult, WriteData,
                input  logic [31:0] ReadData);

  logic [31:0] PCNext, PCPlus4, PCTarget;
  logic [31:0] ImmExt;
  logic [31:0] SrcA, SrcB;
  logic [31:0] Result;

  // next PC logic
  flopr #(32) pcreg(clk, reset, PCNext, PC); // Registrador para o PC
  adder       pcadd4(PC, 32'd4, PCPlus4); // Lógica PC + 4
  adder       pcaddbranch(PC, ImmExt, PCTarget); // Lógica do PC + Imm
  mux2 #(32)  pcmux(PCPlus4, PCTarget, PCSrc, PCNext); // Mux para definir um branch ou fluxo "normal" do PC
 
  // register file logic
  regfile     rf(clk, RegWrite, Instr[19:15], Instr[24:20], 
                 Instr[11:7], Result, SrcA, WriteData);
  extend      ext(Instr[31:7], ImmSrc, ImmExt); // modulo do immediato

  // ALU logic
  mux2 #(32)  srcbmux(WriteData, ImmExt, ALUSrc, SrcB); // Mux para verificar se a soma sera feita com o immediato ou com o rs2
  alu         alu(SrcA, SrcB, ALUControl, ALUResult, Zero); 
  mux3 #(32)  resultmux(ALUResult, ReadData, 32'b0, ResultSrc, Result); // Mux para passar o resultado da ALU direto ou o dado lido da memória
endmodule

// Banco de registradores
module regfile(input  logic        clk, 
               input  logic        we3, 
               input  logic [ 4:0] a1, a2, a3, 
               input  logic [31:0] wd3, 
               output logic [31:0] rd1, rd2);

  logic [31:0] rf[31:0];

  // three ported register file
  // read two ports combinationally (A1/RD1, A2/RD2)
  // write third port on rising edge of clock (A3/WD3/WE3)
  // register 0 hardwired to 0

  always_ff @(posedge clk)
    if (we3) rf[a3] <= wd3;	// Se we3 estiver em alto o dado é escrito no registrador rd(a3)

  assign rd1 = (a1 != 0) ? rf[a1] : 0; // verifica se o registrador rs1(a1) é 0 se for atribui 0 se não a1
  assign rd2 = (a2 != 0) ? rf[a2] : 0; // verifica se o registrador rs20(a2) é 0 se for atribui 0 se não a2
endmodule

// Somador
module adder(input  [31:0] a, b,
             output [31:0] y);

  assign y = a + b;
endmodule

// Modulo Immediato
module extend(input  logic [31:7] instr,
              input  logic [1:0]  immsrc,
              output logic [31:0] immext);
 
  always_comb
    case(immsrc) 
      2'b00:   immext = {{20{instr[31]}}, instr[31:20]};                      // I-type
      2'b01:   immext = {{20{instr[31]}}, instr[31:25], instr[11:7]};         // S-type
      2'b10:   immext = {{20{instr[31]}}, instr[7], instr[30:25], instr[11:8], 1'b0}; // B-type
      2'b11:   immext = {{12{instr[31]}}, instr[19:12], instr[20], instr[30:21], 1'b0}; // J-type
      default: immext = 32'bx; // undefined
    endcase             
endmodule

// Flip Flop genérico
module flopr #(parameter WIDTH = 8)
              (input  logic             clk, reset,
               input  logic [WIDTH-1:0] d, 
               output logic [WIDTH-1:0] q);

  always_ff @(posedge clk, posedge reset)
    if (reset) q <= 0;
    else       q <= d;
endmodule

module mux2 #(parameter WIDTH = 8)
             (input  logic [WIDTH-1:0] d0, d1, 
              input  logic             s, 
              output logic [WIDTH-1:0] y);

  assign y = s ? d1 : d0; 
endmodule

module mux3 #(parameter WIDTH = 8)
             (input  logic [WIDTH-1:0] d0, d1, d2,
              input  logic [1:0]       s, 
              output logic [WIDTH-1:0] y);

  assign y = s[1] ? d2 : (s[0] ? d1 : d0); 
endmodule

module imem(input  logic [31:0] a,
            output logic [31:0] rd);

  logic [31:0] RAM[63:0]; // instancia um array de 64 x 32

  initial
      $readmemh("riscvtest.txt",RAM); // Lê os comandos em hexa baseado em riscv

  assign rd = RAM[a[31:2]]; // word aligned, ou seja acessa a memória 
endmodule

module dmem(input  logic        clk, we,
            input  logic [31:0] a, wd,
            output logic [31:0] rd);

  logic [31:0] RAM[63:0]; // instancia um vetor de memória

  assign rd = RAM[a[31:2]]; // word aligned // atribui a saída rd a o dada da memória e lê o dado se 

  always_ff @(posedge clk) //flip flip de subida do clock
    if (we) RAM[a[31:2]] <= wd; // se o sinal de escrita estiver ativo o valor 
                                // de wd é escrito na memória
endmodule

module alu(input  logic [31:0] a, b,
           input  logic [2:0]  alucontrol,
           output logic [31:0] result,
           output logic        zero);

  logic [31:0] condinvb, sum;
  logic        v;              // overflow
  logic        isAddSub;       // true when is add or subtract operation

  assign condinvb = alucontrol[0] ? ~b : b;
  assign sum = a + condinvb + alucontrol[0];
  assign isAddSub = ~alucontrol[2] & ~alucontrol[1] |
                    ~alucontrol[1] & alucontrol[0];

  always_comb
    case (alucontrol)
      3'b000:  result = sum;         // add
      3'b001:  result = sum;         // subtract
      3'b010:  result = a & b;       // and
      3'b011:  result = a | b;       // or
      3'b100:  result = a ^ b;       // xor
      3'b101:  result = sum[31] ^ v; // slt
      3'b110:  result = a << b[4:0]; // sll
      3'b111:  result = a >> b[4:0]; // srl
      default: result = 32'bx;
    endcase

  assign zero = (result == 32'b0);
  assign v = ~(alucontrol[0] ^ a[31] ^ b[31]) & (a[31] ^ sum[31]) & isAddSub;
  
endmodule
